.subckt opamp vinp vinn vout vdd gnd
m1      d1    vinp  s1  vdd pmos_3p3 L='l_fixed*1u' W='w1_2*1u'
m2      d2    vinn  s1  vdd pmos_3p3 L='l_fixed*1u' W='w1_2*1u'
m3      d3    vinp  s3  gnd nmos_3p3 L='l_fixed*1u' W='w3_4*1u'
m4      d4    vinn  s3  gnd nmos_3p3 L='l_fixed*1u' W='w3_4*1u'
m5      s1    g5    vdd vdd pmos_3p3 L='l_fixed*1u' w='w5*1u'
m6      s3    ibias gnd gnd nmos_3p3 L='l_fixed*1u' w='w6*1u'
m7      ibias ibias gnd gnd nmos_3p3 L='l_fixed*1u' w='w7*1u'
m8      g5    ibias gnd gnd nmos_3p3 L='l_fixed*1u' w='w8*1u'
m9      g5    g5    vdd vdd pmos_3p3 L='l_fixed*1u' w='w9*1u'
m10     d10   ibias gnd gnd nmos_3p3 L='l_fixed*1u' w='w10*1u'
m11     d10   d10   s11 vdd pmos_3p3 L='l_fixed*1u' w='w11*1u'
m12     s11   d10   vdd vdd pmos_3p3 L='l_fixed*1u' w='w12*1u'
m13     d13   g5    vdd vdd pmos_3p3 L='l_fixed*1u' w='w13*1u'
m14     d13   d13   s14 gnd nmos_3p3 L='l_fixed*1u' w='w14*1u'
m15     s14   d13   gnd gnd nmos_3p3 L='l_fixed*1u' w='w15*1u'
m16     d16   d13   d2  gnd nmos_3p3 L='l_fixed*1u' W='w16_18*1u'
m17     d2    d16   gnd gnd nmos_3p3 L='l_fixed*1u' W='w17_19*1u'
m18     d18   d13   d1  gnd nmos_3p3 L='l_fixed*1u' W='w16_18*1u'
m19     d1    d16   gnd gnd nmos_3p3 L='l_fixed*1u' W='w17_19*1u'
m20     d16   d10   d4  vdd pmos_3p3 L='l_fixed*1u' W='w20*1u'
m21     d21   d10   d3  vdd pmos_3p3 L='l_fixed*1u' W='w21*1u'
m22     d4    g5    vdd vdd pmos_3p3 L='l_fixed*1u' W='w22_23*1u'
m23     d3    g5    vdd vdd pmos_3p3 L='l_fixed*1u' W='w22_23*1u'
m24     d24   g5    vdd vdd pmos_3p3 L='l_fixed*1u' W='w24*1u'
m25     d25   d10   d24 vdd pmos_3p3 L='l_fixed*1u' W='w25*1u'
m26     d25   d25   s26 gnd nmos_3p3 L='l_fixed*1u' W='w26*1u'
m27     s26   s26   gnd gnd nmos_3p3 L='l_fixed*1u' W='w27*1u'
m28     d28   ibias gnd gnd nmos_3p3 L='l_fixed*1u' W='w28*1u'
m29     d29   d13   d28 gnd nmos_3p3 L='l_fixed*1u' W='w29*1u'
m30     d29   d29   s30 vdd pmos_3p3 L='l_fixed*1u' W='w30*1u'
m31     s30   s30   vdd vdd pmos_3p3 L='l_fixed*1u' W='w31*1u'
m32     vout  d21   vdd vdd pmos_3p3 L='l_fixed*1u' W='w32*1u'
m33     vout  d18   gnd gnd nmos_3p3 L='l_fixed*1u' W='w33*1u'
m34     d21   d25   d18 gnd nmos_3p3 L='l_fixed*1u' W='w34*1u'
m35     d18   d29   d21 vdd pmos_3p3 L='l_fixed*1u' w='w35*1u'
ibias vdd ibias dc='ival*1e-3'
cm d1 vout 'cm*1p'
cload vout gnd 1p 
.ENDS
