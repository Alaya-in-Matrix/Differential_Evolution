.if(weff1_2 > 20)
.param m1_2 = 2
.else
.param m1_2 = 1
.endif
.if(weff3_4 > 20)
.param m3_4 = 2
.else
.param m3_4 = 1
.endif
.if(weff5 > 20)
.param m5 = 2
.else
.param m5 = 1
.endif
.if(weff6 > 20)
.param m6 = 2
.else
.param m6 = 1
.endif
.if(weff7 > 20)
.param m7 = 2
.else
.param m7 = 1
.endif
.if(weff8 > 20)
.param m8 = 2
.else
.param m8 = 1
.endif
.if(weff9 > 20)
.param m9 = 2
.else
.param m9 = 1
.endif
.if(weff10 > 20)
.param m10 = 2
.else
.param m10 = 1
.endif
.if(weff11 > 20)
.param m11 = 2
.else
.param m11 = 1
.endif
.if(weff12 > 20)
.param m12 = 2
.else
.param m12 = 1
.endif
.if(weff13 > 20)
.param m13 = 2
.else
.param m13 = 1
.endif
.if(weff14 > 20)
.param m14 = 2
.else
.param m14 = 1
.endif
.if(weff15 > 20)
.param m15 = 2
.else
.param m15 = 1
.endif
.if(weff16_18 > 20)
.param m16_18 = 2
.else
.param m16_18 = 1
.endif
.if(weff17_19 > 20)
.param m17_19 = 2
.else
.param m17_19 = 1
.endif
.if(weff20 > 20)
.param m20 = 2
.else
.param m20 = 1
.endif
.if(weff21 > 20)
.param m21 = 2
.else
.param m21 = 1
.endif
.if(weff22_23 > 20)
.param m22_23 = 2
.else
.param m22_23 = 1
.endif
.if(weff24 > 20)
.param m24 = 2
.else
.param m24 = 1
.endif
.if(weff25 > 20)
.param m25 = 2
.else
.param m25 = 1
.endif
.if(weff26 > 20)
.param m26 = 2
.else
.param m26 = 1
.endif
.if(weff27 > 20)
.param m27 = 2
.else
.param m27 = 1
.endif
.if(weff28 > 20)
.param m28 = 2
.else
.param m28 = 1
.endif
.if(weff29 > 20)
.param m29 = 2
.else
.param m29 = 1
.endif
.if(weff30 > 20)
.param m30 = 2
.else
.param m30 = 1
.endif
.if(weff31 > 20)
.param m31 = 2
.else
.param m31 = 1
.endif
.if(weff32 > 20)
.param m32 = 2
.else
.param m32 = 1
.endif
.if(weff33 > 20)
.param m33 = 2
.else
.param m33 = 1
.endif
.if(weff34 > 20)
.param m34 = 2
.else
.param m34 = 1
.endif
.if(weff35 > 20)
.param m35 = 2
.else
.param m35 = 1
.endif
.param w1_2   = 'weff1_2/m1_2'
.param w3_4   = 'weff3_4/m3_4'
.param w5     = 'weff5/m5'
.param w6     = 'weff6/m6'
.param w7     = 'weff7/m7'
.param w8     = 'weff8/m8'
.param w9     = 'weff9/m9'
.param w10    = 'weff10/m10'
.param w11    = 'weff11/m11'
.param w12    = 'weff12/m12'
.param w13    = 'weff13/m13'
.param w14    = 'weff14/m14'
.param w15    = 'weff15/m15'
.param w16_18 = 'weff16_18/m16_18'
.param w17_19 = 'weff17_19/m17_19'
.param w20    = 'weff20/m20'
.param w21    = 'weff21/m21'
.param w22_23 = 'weff22_23/m22_23'
.param w24    = 'weff24/m24'
.param w25    = 'weff25/m25'
.param w26    = 'weff26/m26'
.param w27    = 'weff27/m27'
.param w28    = 'weff28/m28'
.param w29    = 'weff29/m29'
.param w30    = 'weff30/m30'
.param w31    = 'weff31/m31'
.param w32    = 'weff32/m32'
.param w33    = 'weff33/m33'
.param w34    = 'weff34/m34'
.param w35    = 'weff35/m35'
